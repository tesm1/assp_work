package myProssu_params is
  constant fu_stream_out_statusw : integer := 8;
  constant fu_stream_in_statusw : integer := 8;
  constant fu_LSU_dataw : integer := 32;
  constant fu_LSU_addrw : integer := 8;
end myProssu_params;
