package myProssu_imem_mau is
   -- created by generatebits
   constant IMEMMAUWIDTH : positive := 344;
end myProssu_imem_mau;
